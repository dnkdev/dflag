module dflag

fn test_parse_struct() {
}
